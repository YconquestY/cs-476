`timescale 1ps/1ps

module wrTxTb;
endmodule