`timescale 1ps/1ps

module rdErrTb;
endmodule